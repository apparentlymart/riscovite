module cpu();

endmodule
